** Profile: "SCHEMATIC1-1"  [ C:\Users\21116132\Documents\Elec_Analog\TP5_PARTIE1-2\tp51-SCHEMATIC1-1.sim ] 

** Creating circuit file "tp51-SCHEMATIC1-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 20 1Hz 1MEGHz
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tp51-SCHEMATIC1.net" 


.END
