** Profile: "SCHEMATIC1-2.2"  [ C:\Users\21116132\Documents\Elec_Analog\TP5_PARTIE1-2\tp51-SCHEMATIC1-2.2.sim ] 

** Creating circuit file "tp51-SCHEMATIC1-2.2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 20 1Hz 1MEGHz
.STEP PARAM val LIST 79.57,7.957k,79.57k,795.774k 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tp51-SCHEMATIC1.net" 


.END
